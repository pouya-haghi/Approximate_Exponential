library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMfact is
    Port ( add : in  STD_LOGIC_VECTOR (3 downto 0);
           data : out  STD_LOGIC_VECTOR (31 downto 0));
end ROMfact;

architecture Behavioral of ROMfact is
begin
with add select
data<=(others=>'1') when "0000",
      "10000000000000000000000000000000" when "0001",
	  "01010101010101010101010101010101" when "0010",
	  "01000000000000000000000000000000" when "0011",
	  "00110011001100110011001100110011" when "0100",
	  "00101010101010101010101010101010" when "0101",
	  "00100100100100100100100100100100" when "0110",
	  "00100000000000000000000000000000" when "0111",
	  "00011100011100011100011100011100" when "1000",
      "00011001100110011001100110011001" when "1001",
	  "00010111010001011101000101110100" when "1010",
	  "00010101010101010101010101010101" when "1011",
	  "00010011101100010011101100010011" when "1100",
	  "00010010010010010010010010010010" when "1101",
	  "00010001000100010001000100010001" when "1110",
	  "00010000000000000000000000000000" when "1111",
	  (others=>'1') when others;
end Behavioral;

